`ifndef MAC_DEFINE_SVH
`define MAC_DEFINE_SVH

// MAC / Ethernet Frame Sizes
`define DST_MAC_BYTES   6
`define SRC_MAC_BYTES   6
`define VLAN_ID_BITS    12
`define PCP_BITS        3
`define DEI_BITS        1
`define ETH_TYPE_BYTES  2
`define MIN_PAYLOAD     46
`define MAX_PAYLOAD     1500
`define FCS_BYTES       4

`endif // MAC_DEFINE_SVH

