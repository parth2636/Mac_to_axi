/* -.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.

* File Name : c2n_mac_lyr_sequencer.sv

* Purpose :

* Creation Date : 13-05-2024

* Last Modified :

* Created By :  

_._._._._._._._._._._._._._._._._._._._._.*/


`ifndef C2N_MAC_LYR_SEQUENCER_SV
`define C2N_MAC_LYR_SEQUENCER_SV

class c2n_mac_lyr_sequencer extends uvm_sequencer; 
 
  `uvm_component_utils(c2n_mac_lyr_sequencer) 
   
    //-------------------------------------------------------------------------------- 
     // Method : 
      
       // Arguments : 
        
         // Description : 
          
           //--------------------------------------------------------------------------------- 
             function new (string name="c2n_mac_lyr_sequencer", uvm_component parent=null); 
               super.new(name,parent); 
                
                  endfunction: new 
                   
                    
                     
                      
                       
                        
                         
                          
                           endclass : c2n_mac_lyr_sequencer


`endif
